`timescale 1ns/1ns

package yapp_pkg;
  import uvm_pkg::*;
  //declaration 
  typedef uvm_config_db#(virtual yapp_if) yapp_vif_config;

  `include "uvm_macros.svh"
  
  `include "../tb/yapp_packet.sv"
  `include "../tb/yapp_tx_monitor.sv"
  `include "../tb/yapp_tx_sequencer.sv"
  `include "../tb/yapp_tx_seqs.sv"
  `include "../tb/yapp_tx_driver.sv"
  `include "../tb/yapp_tx_agent.sv"
  `include "../tb/yapp_tx_env.sv"
  
endpackage